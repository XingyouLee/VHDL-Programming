--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   09:19:58 05/14/2021
-- Design Name:   
-- Module Name:   C:/Users/XingyouLee/OneDrive/Program/VHDL/test1/atest.vhd
-- Project Name:  test1
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: test1
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY atest IS
END atest;
 
ARCHITECTURE behavior OF atest IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT test1
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         taken : IN  std_logic;
         predict : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';
   signal taken : std_logic := '0';

 	--Outputs
   signal predict : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: test1 PORT MAP (
          clk => clk,
          reset => reset,
          taken => taken,
          predict => predict
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      reset <= '1';
      wait for 10 ns;
      taken <= '0';
      wait for 100 ns;
      taken <= '0';
      wait for 100 ns;
      taken <= '0';
      wait for 100 ns;
      taken <= '1';
      wait for 100 ns;
      taken <= '1';
      wait for 100 ns;

      wait;
   end process;

END;
